module helpers

pub fn blue() string {
	return '\e[0;34m'
}

pub fn reset() string {
	return '\e[0m'
}